// system.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module system (
		input  wire        ad9276_spi_external_MISO,       //     ad9276_spi_external.MISO
		output wire        ad9276_spi_external_MOSI,       //                        .MOSI
		output wire        ad9276_spi_external_SCLK,       //                        .SCLK
		output wire        ad9276_spi_external_SS_n,       //                        .SS_n
		input  wire        clk_clk,                        //                     clk.clk
		input  wire [69:0] datain_probe,                   //                  datain.probe
		output wire [69:0] dataout_source,                 //                 dataout.source
		output wire [31:0] general_cnt_export,             //             general_cnt.export
		output wire [9:0]  issp_cnt_source,                //                issp_cnt.source
		output wire [31:0] lm96570_spi_in_0_export,        //        lm96570_spi_in_0.export
		output wire [31:0] lm96570_spi_in_1_export,        //        lm96570_spi_in_1.export
		output wire [5:0]  lm96570_spi_in_2_export,        //        lm96570_spi_in_2.export
		output wire [7:0]  lm96570_spi_num_of_bits_export, // lm96570_spi_num_of_bits.export
		input  wire [31:0] lm96570_spi_out_0_export,       //       lm96570_spi_out_0.export
		input  wire [31:0] lm96570_spi_out_1_export,       //       lm96570_spi_out_1.export
		input  wire [5:0]  lm96570_spi_out_2_export,       //       lm96570_spi_out_2.export
		output wire [7:0]  num_of_bits_source,             //             num_of_bits.source
		output wire        pll_0_locked_export,            //            pll_0_locked.export
		output wire        pll_0_outclk0_clk,              //           pll_0_outclk0.clk
		input  wire        reset_reset_n                   //                   reset.reset_n
	);

	wire  [31:0] master_0_master_readdata;                                 // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                              // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                  // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                     // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                               // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                            // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                    // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire         mm_interconnect_0_lm96570_spi_in_2_s1_chipselect;         // mm_interconnect_0:lm96570_spi_in_2_s1_chipselect -> lm96570_spi_in_2:chipselect
	wire  [31:0] mm_interconnect_0_lm96570_spi_in_2_s1_readdata;           // lm96570_spi_in_2:readdata -> mm_interconnect_0:lm96570_spi_in_2_s1_readdata
	wire   [1:0] mm_interconnect_0_lm96570_spi_in_2_s1_address;            // mm_interconnect_0:lm96570_spi_in_2_s1_address -> lm96570_spi_in_2:address
	wire         mm_interconnect_0_lm96570_spi_in_2_s1_write;              // mm_interconnect_0:lm96570_spi_in_2_s1_write -> lm96570_spi_in_2:write_n
	wire  [31:0] mm_interconnect_0_lm96570_spi_in_2_s1_writedata;          // mm_interconnect_0:lm96570_spi_in_2_s1_writedata -> lm96570_spi_in_2:writedata
	wire         mm_interconnect_0_lm96570_spi_in_0_s1_chipselect;         // mm_interconnect_0:lm96570_spi_in_0_s1_chipselect -> lm96570_spi_in_0:chipselect
	wire  [31:0] mm_interconnect_0_lm96570_spi_in_0_s1_readdata;           // lm96570_spi_in_0:readdata -> mm_interconnect_0:lm96570_spi_in_0_s1_readdata
	wire   [1:0] mm_interconnect_0_lm96570_spi_in_0_s1_address;            // mm_interconnect_0:lm96570_spi_in_0_s1_address -> lm96570_spi_in_0:address
	wire         mm_interconnect_0_lm96570_spi_in_0_s1_write;              // mm_interconnect_0:lm96570_spi_in_0_s1_write -> lm96570_spi_in_0:write_n
	wire  [31:0] mm_interconnect_0_lm96570_spi_in_0_s1_writedata;          // mm_interconnect_0:lm96570_spi_in_0_s1_writedata -> lm96570_spi_in_0:writedata
	wire         mm_interconnect_0_lm96570_spi_in_1_s1_chipselect;         // mm_interconnect_0:lm96570_spi_in_1_s1_chipselect -> lm96570_spi_in_1:chipselect
	wire  [31:0] mm_interconnect_0_lm96570_spi_in_1_s1_readdata;           // lm96570_spi_in_1:readdata -> mm_interconnect_0:lm96570_spi_in_1_s1_readdata
	wire   [1:0] mm_interconnect_0_lm96570_spi_in_1_s1_address;            // mm_interconnect_0:lm96570_spi_in_1_s1_address -> lm96570_spi_in_1:address
	wire         mm_interconnect_0_lm96570_spi_in_1_s1_write;              // mm_interconnect_0:lm96570_spi_in_1_s1_write -> lm96570_spi_in_1:write_n
	wire  [31:0] mm_interconnect_0_lm96570_spi_in_1_s1_writedata;          // mm_interconnect_0:lm96570_spi_in_1_s1_writedata -> lm96570_spi_in_1:writedata
	wire  [31:0] mm_interconnect_0_lm96570_spi_out_2_s1_readdata;          // lm96570_spi_out_2:readdata -> mm_interconnect_0:lm96570_spi_out_2_s1_readdata
	wire   [1:0] mm_interconnect_0_lm96570_spi_out_2_s1_address;           // mm_interconnect_0:lm96570_spi_out_2_s1_address -> lm96570_spi_out_2:address
	wire  [31:0] mm_interconnect_0_lm96570_spi_out_1_s1_readdata;          // lm96570_spi_out_1:readdata -> mm_interconnect_0:lm96570_spi_out_1_s1_readdata
	wire   [1:0] mm_interconnect_0_lm96570_spi_out_1_s1_address;           // mm_interconnect_0:lm96570_spi_out_1_s1_address -> lm96570_spi_out_1:address
	wire  [31:0] mm_interconnect_0_lm96570_spi_out_0_s1_readdata;          // lm96570_spi_out_0:readdata -> mm_interconnect_0:lm96570_spi_out_0_s1_readdata
	wire   [1:0] mm_interconnect_0_lm96570_spi_out_0_s1_address;           // mm_interconnect_0:lm96570_spi_out_0_s1_address -> lm96570_spi_out_0:address
	wire         mm_interconnect_0_lm96570_spi_num_of_bits_s1_chipselect;  // mm_interconnect_0:lm96570_spi_num_of_bits_s1_chipselect -> lm96570_spi_num_of_bits:chipselect
	wire  [31:0] mm_interconnect_0_lm96570_spi_num_of_bits_s1_readdata;    // lm96570_spi_num_of_bits:readdata -> mm_interconnect_0:lm96570_spi_num_of_bits_s1_readdata
	wire   [1:0] mm_interconnect_0_lm96570_spi_num_of_bits_s1_address;     // mm_interconnect_0:lm96570_spi_num_of_bits_s1_address -> lm96570_spi_num_of_bits:address
	wire         mm_interconnect_0_lm96570_spi_num_of_bits_s1_write;       // mm_interconnect_0:lm96570_spi_num_of_bits_s1_write -> lm96570_spi_num_of_bits:write_n
	wire  [31:0] mm_interconnect_0_lm96570_spi_num_of_bits_s1_writedata;   // mm_interconnect_0:lm96570_spi_num_of_bits_s1_writedata -> lm96570_spi_num_of_bits:writedata
	wire         mm_interconnect_0_general_cnt_s1_chipselect;              // mm_interconnect_0:general_cnt_s1_chipselect -> general_cnt:chipselect
	wire  [31:0] mm_interconnect_0_general_cnt_s1_readdata;                // general_cnt:readdata -> mm_interconnect_0:general_cnt_s1_readdata
	wire   [1:0] mm_interconnect_0_general_cnt_s1_address;                 // mm_interconnect_0:general_cnt_s1_address -> general_cnt:address
	wire         mm_interconnect_0_general_cnt_s1_write;                   // mm_interconnect_0:general_cnt_s1_write -> general_cnt:write_n
	wire  [31:0] mm_interconnect_0_general_cnt_s1_writedata;               // mm_interconnect_0:general_cnt_s1_writedata -> general_cnt:writedata
	wire         mm_interconnect_0_ad9276_spi_spi_control_port_chipselect; // mm_interconnect_0:ad9276_spi_spi_control_port_chipselect -> ad9276_spi:spi_select
	wire  [31:0] mm_interconnect_0_ad9276_spi_spi_control_port_readdata;   // ad9276_spi:data_to_cpu -> mm_interconnect_0:ad9276_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_ad9276_spi_spi_control_port_address;    // mm_interconnect_0:ad9276_spi_spi_control_port_address -> ad9276_spi:mem_addr
	wire         mm_interconnect_0_ad9276_spi_spi_control_port_read;       // mm_interconnect_0:ad9276_spi_spi_control_port_read -> ad9276_spi:read_n
	wire         mm_interconnect_0_ad9276_spi_spi_control_port_write;      // mm_interconnect_0:ad9276_spi_spi_control_port_write -> ad9276_spi:write_n
	wire  [31:0] mm_interconnect_0_ad9276_spi_spi_control_port_writedata;  // mm_interconnect_0:ad9276_spi_spi_control_port_writedata -> ad9276_spi:data_from_cpu
	wire         rst_controller_reset_out_reset;                           // rst_controller:reset_out -> [ad9276_spi:reset_n, general_cnt:reset_n, lm96570_spi_in_0:reset_n, lm96570_spi_in_1:reset_n, lm96570_spi_in_2:reset_n, lm96570_spi_num_of_bits:reset_n, lm96570_spi_out_0:reset_n, lm96570_spi_out_1:reset_n, lm96570_spi_out_2:reset_n, mm_interconnect_0:lm96570_spi_in_2_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset]

	system_ad9276_spi ad9276_spi (
		.clk           (clk_clk),                                                  //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                          //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_ad9276_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_ad9276_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_ad9276_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_ad9276_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_ad9276_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_ad9276_spi_spi_control_port_write),     //                 .write_n
		.irq           (),                                                         //              irq.irq
		.MISO          (ad9276_spi_external_MISO),                                 //         external.export
		.MOSI          (ad9276_spi_external_MOSI),                                 //                 .export
		.SCLK          (ad9276_spi_external_SCLK),                                 //                 .export
		.SS_n          (ad9276_spi_external_SS_n)                                  //                 .export
	);

	system_general_cnt general_cnt (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_general_cnt_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_general_cnt_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_general_cnt_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_general_cnt_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_general_cnt_s1_readdata),   //                    .readdata
		.out_port   (general_cnt_export)                           // external_connection.export
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("NONE"),
		.probe_width             (70),
		.source_width            (70),
		.source_initial_value    ("0"),
		.enable_metastability    ("NO")
	) in_system_sources_probes_0 (
		.source     (dataout_source), // sources.source
		.probe      (datain_probe),   //  probes.probe
		.source_ena (1'b1)            // (terminated)
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("NONE"),
		.probe_width             (0),
		.source_width            (8),
		.source_initial_value    ("0"),
		.enable_metastability    ("NO")
	) in_system_sources_probes_1 (
		.source     (num_of_bits_source), // sources.source
		.source_ena (1'b1)                // (terminated)
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("NONE"),
		.probe_width             (0),
		.source_width            (10),
		.source_initial_value    ("0"),
		.enable_metastability    ("NO")
	) in_system_sources_probes_2 (
		.source     (issp_cnt_source), // sources.source
		.source_ena (1'b1)             // (terminated)
	);

	system_general_cnt lm96570_spi_in_0 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_lm96570_spi_in_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lm96570_spi_in_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lm96570_spi_in_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lm96570_spi_in_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lm96570_spi_in_0_s1_readdata),   //                    .readdata
		.out_port   (lm96570_spi_in_0_export)                           // external_connection.export
	);

	system_general_cnt lm96570_spi_in_1 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_lm96570_spi_in_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lm96570_spi_in_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lm96570_spi_in_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lm96570_spi_in_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lm96570_spi_in_1_s1_readdata),   //                    .readdata
		.out_port   (lm96570_spi_in_1_export)                           // external_connection.export
	);

	system_lm96570_spi_in_2 lm96570_spi_in_2 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_lm96570_spi_in_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lm96570_spi_in_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lm96570_spi_in_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lm96570_spi_in_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lm96570_spi_in_2_s1_readdata),   //                    .readdata
		.out_port   (lm96570_spi_in_2_export)                           // external_connection.export
	);

	system_lm96570_spi_num_of_bits lm96570_spi_num_of_bits (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (mm_interconnect_0_lm96570_spi_num_of_bits_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lm96570_spi_num_of_bits_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lm96570_spi_num_of_bits_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lm96570_spi_num_of_bits_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lm96570_spi_num_of_bits_s1_readdata),   //                    .readdata
		.out_port   (lm96570_spi_num_of_bits_export)                           // external_connection.export
	);

	system_lm96570_spi_out_0 lm96570_spi_out_0 (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_lm96570_spi_out_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_lm96570_spi_out_0_s1_readdata), //                    .readdata
		.in_port  (lm96570_spi_out_0_export)                         // external_connection.export
	);

	system_lm96570_spi_out_0 lm96570_spi_out_1 (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_lm96570_spi_out_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_lm96570_spi_out_1_s1_readdata), //                    .readdata
		.in_port  (lm96570_spi_out_1_export)                         // external_connection.export
	);

	system_lm96570_spi_out_2 lm96570_spi_out_2 (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_lm96570_spi_out_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_lm96570_spi_out_2_s1_readdata), //                    .readdata
		.in_port  (lm96570_spi_out_2_export)                         // external_connection.export
	);

	system_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	system_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),   // outclk0.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                      (clk_clk),                                                  //                                    clk_0_clk.clk
		.lm96570_spi_in_2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                           // lm96570_spi_in_2_reset_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                           //     master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_address                            (master_0_master_address),                                  //                              master_0_master.address
		.master_0_master_waitrequest                        (master_0_master_waitrequest),                              //                                             .waitrequest
		.master_0_master_byteenable                         (master_0_master_byteenable),                               //                                             .byteenable
		.master_0_master_read                               (master_0_master_read),                                     //                                             .read
		.master_0_master_readdata                           (master_0_master_readdata),                                 //                                             .readdata
		.master_0_master_readdatavalid                      (master_0_master_readdatavalid),                            //                                             .readdatavalid
		.master_0_master_write                              (master_0_master_write),                                    //                                             .write
		.master_0_master_writedata                          (master_0_master_writedata),                                //                                             .writedata
		.ad9276_spi_spi_control_port_address                (mm_interconnect_0_ad9276_spi_spi_control_port_address),    //                  ad9276_spi_spi_control_port.address
		.ad9276_spi_spi_control_port_write                  (mm_interconnect_0_ad9276_spi_spi_control_port_write),      //                                             .write
		.ad9276_spi_spi_control_port_read                   (mm_interconnect_0_ad9276_spi_spi_control_port_read),       //                                             .read
		.ad9276_spi_spi_control_port_readdata               (mm_interconnect_0_ad9276_spi_spi_control_port_readdata),   //                                             .readdata
		.ad9276_spi_spi_control_port_writedata              (mm_interconnect_0_ad9276_spi_spi_control_port_writedata),  //                                             .writedata
		.ad9276_spi_spi_control_port_chipselect             (mm_interconnect_0_ad9276_spi_spi_control_port_chipselect), //                                             .chipselect
		.general_cnt_s1_address                             (mm_interconnect_0_general_cnt_s1_address),                 //                               general_cnt_s1.address
		.general_cnt_s1_write                               (mm_interconnect_0_general_cnt_s1_write),                   //                                             .write
		.general_cnt_s1_readdata                            (mm_interconnect_0_general_cnt_s1_readdata),                //                                             .readdata
		.general_cnt_s1_writedata                           (mm_interconnect_0_general_cnt_s1_writedata),               //                                             .writedata
		.general_cnt_s1_chipselect                          (mm_interconnect_0_general_cnt_s1_chipselect),              //                                             .chipselect
		.lm96570_spi_in_0_s1_address                        (mm_interconnect_0_lm96570_spi_in_0_s1_address),            //                          lm96570_spi_in_0_s1.address
		.lm96570_spi_in_0_s1_write                          (mm_interconnect_0_lm96570_spi_in_0_s1_write),              //                                             .write
		.lm96570_spi_in_0_s1_readdata                       (mm_interconnect_0_lm96570_spi_in_0_s1_readdata),           //                                             .readdata
		.lm96570_spi_in_0_s1_writedata                      (mm_interconnect_0_lm96570_spi_in_0_s1_writedata),          //                                             .writedata
		.lm96570_spi_in_0_s1_chipselect                     (mm_interconnect_0_lm96570_spi_in_0_s1_chipselect),         //                                             .chipselect
		.lm96570_spi_in_1_s1_address                        (mm_interconnect_0_lm96570_spi_in_1_s1_address),            //                          lm96570_spi_in_1_s1.address
		.lm96570_spi_in_1_s1_write                          (mm_interconnect_0_lm96570_spi_in_1_s1_write),              //                                             .write
		.lm96570_spi_in_1_s1_readdata                       (mm_interconnect_0_lm96570_spi_in_1_s1_readdata),           //                                             .readdata
		.lm96570_spi_in_1_s1_writedata                      (mm_interconnect_0_lm96570_spi_in_1_s1_writedata),          //                                             .writedata
		.lm96570_spi_in_1_s1_chipselect                     (mm_interconnect_0_lm96570_spi_in_1_s1_chipselect),         //                                             .chipselect
		.lm96570_spi_in_2_s1_address                        (mm_interconnect_0_lm96570_spi_in_2_s1_address),            //                          lm96570_spi_in_2_s1.address
		.lm96570_spi_in_2_s1_write                          (mm_interconnect_0_lm96570_spi_in_2_s1_write),              //                                             .write
		.lm96570_spi_in_2_s1_readdata                       (mm_interconnect_0_lm96570_spi_in_2_s1_readdata),           //                                             .readdata
		.lm96570_spi_in_2_s1_writedata                      (mm_interconnect_0_lm96570_spi_in_2_s1_writedata),          //                                             .writedata
		.lm96570_spi_in_2_s1_chipselect                     (mm_interconnect_0_lm96570_spi_in_2_s1_chipselect),         //                                             .chipselect
		.lm96570_spi_num_of_bits_s1_address                 (mm_interconnect_0_lm96570_spi_num_of_bits_s1_address),     //                   lm96570_spi_num_of_bits_s1.address
		.lm96570_spi_num_of_bits_s1_write                   (mm_interconnect_0_lm96570_spi_num_of_bits_s1_write),       //                                             .write
		.lm96570_spi_num_of_bits_s1_readdata                (mm_interconnect_0_lm96570_spi_num_of_bits_s1_readdata),    //                                             .readdata
		.lm96570_spi_num_of_bits_s1_writedata               (mm_interconnect_0_lm96570_spi_num_of_bits_s1_writedata),   //                                             .writedata
		.lm96570_spi_num_of_bits_s1_chipselect              (mm_interconnect_0_lm96570_spi_num_of_bits_s1_chipselect),  //                                             .chipselect
		.lm96570_spi_out_0_s1_address                       (mm_interconnect_0_lm96570_spi_out_0_s1_address),           //                         lm96570_spi_out_0_s1.address
		.lm96570_spi_out_0_s1_readdata                      (mm_interconnect_0_lm96570_spi_out_0_s1_readdata),          //                                             .readdata
		.lm96570_spi_out_1_s1_address                       (mm_interconnect_0_lm96570_spi_out_1_s1_address),           //                         lm96570_spi_out_1_s1.address
		.lm96570_spi_out_1_s1_readdata                      (mm_interconnect_0_lm96570_spi_out_1_s1_readdata),          //                                             .readdata
		.lm96570_spi_out_2_s1_address                       (mm_interconnect_0_lm96570_spi_out_2_s1_address),           //                         lm96570_spi_out_2_s1.address
		.lm96570_spi_out_2_s1_readdata                      (mm_interconnect_0_lm96570_spi_out_2_s1_readdata)           //                                             .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
